
// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   CPU.rf
`define DMEM_PATH CPU.dmem
`define IMEM_PATH CPU.imem

