
// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   CPU.id.rf
`define DMEM_PATH CPU.ex.dmem
`define IMEM_PATH CPU.imem

